-- $File: LED.vhd
-- $Date: Wed Mar 13 20:52:51 2013 +0800
-- $Author: jiakai <jia.kai66@gmail.com>
